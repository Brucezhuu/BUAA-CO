`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:57:05 12/08/2021 
// Design Name: 
// Module Name:    test_shift 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module test_shift(
    input [31:0] rs,
    input [31:0] rt,
    input [31:0] rd,
    output [31:0] res
    );
	
	
	
endmodule
